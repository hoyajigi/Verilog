`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:19:13 03/12/2013 
// Design Name: 
// Module Name:    CA_Inv 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module CA_Inv(In,Out
    );
	input In;
	output Out;
	wire Out;
	
	assign Out=~In;


endmodule
