----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:48:33 06/05/2013 
-- Design Name: 
-- Module Name:    MIPS_Datapath - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MIPS_Datapath is
    Port ( clk : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           TestPort : out  STD_LOGIC_VECTOR (31 downto 0));
end MIPS_Datapath;

architecture Behavioral of MIPS_Datapath is

begin


end Behavioral;

