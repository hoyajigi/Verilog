`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:57:00 03/12/2013 
// Design Name: 
// Module Name:    CA_AND2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module CA_AND2(In1,In2,Out
    );
	input In1,In2;
	output Out;
	wire Out;
	
	assign Out = In1& In2;

endmodule
